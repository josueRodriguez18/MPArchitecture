module riscCPU()